`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09.12.2020 23:21:20
// Design Name: 
// Module Name: snaketop
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



`timescale 1ns/1ps
module alpha1(hpos, vpos, alpha_s);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_s;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-100;
  wire [9:0] y = vpos-200;
  
  assign alpha_s= ((100<=hpos)&(hpos<=149))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
    maze[0]  = 50'b11111111111111111111111111111111111111111111111111; 
 	maze[1]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[2]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[3]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[4]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[5]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[6]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[7]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[8]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[9]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[10] = 50'b11111111111100000000000000000000000000000000000000;
    maze[11] = 50'b11111111111100000000000000000000000000000000000000;
    maze[12] = 50'b11111111111100000000000000000000000000000000000000;
    maze[13] = 50'b11111111111100000000000000000000000000000000000000;
    maze[14] = 50'b11111111111100000000000000000000000000000000000000;
    maze[15] = 50'b11111111111100000000000000000000000000000000000000;
    maze[16] = 50'b11111111111100000000000000000000000000000000000000;
    maze[17] = 50'b11111111111100000000000000000000000000000000000000;
    maze[18] = 50'b11111111111100000000000000000000000000000000000000;
    maze[19] = 50'b11111111111100000000000000000000000000000000000000;
    maze[20] = 50'b11111111111100000000000000000000000000000000000000;
    maze[21] = 50'b11111111111100000000000000000000000000000000000000;
    maze[22] = 50'b11111111111100000000000000000000000000000000000000;
    maze[23] = 50'b11111111111111111111111111111111111111111111111111;
    maze[24] = 50'b11111111111111111111111111111111111111111111111111;
    maze[25] = 50'b11111111111111111111111111111111111111111111111111;
    maze[26] = 50'b11111111111111111111111111111111111111111111111111;
    maze[27] = 50'b11111111111111111111111111111111111111111111111111;
    maze[28] = 50'b00000000000000000000000000000000000000111111111111;
    maze[29] = 50'b00000000000000000000000000000000000000111111111111;
    maze[30] = 50'b00000000000000000000000000000000000000111111111111;
    maze[31] = 50'b00000000000000000000000000000000000000111111111111;
    maze[32] = 50'b00000000000000000000000000000000000000111111111111;
    maze[33] = 50'b00000000000000000000000000000000000000111111111111;
    maze[34] = 50'b00000000000000000000000000000000000000111111111111;
    maze[35] = 50'b00000000000000000000000000000000000000111111111111;
    maze[36] = 50'b00000000000000000000000000000000000000111111111111;
    maze[37] = 50'b00000000000000000000000000000000000000111111111111;
    maze[38] = 50'b00000000000000000000000000000000000000111111111111;
    maze[39] = 50'b00000000000000000000000000000000000000111111111111;
    maze[40] = 50'b00000000000000000000000000000000000000111111111111;
    maze[41] = 50'b00000000000000000000000000000000000000111111111111;
    maze[42] = 50'b00000000000000000000000000000000000000111111111111;
    maze[43] = 50'b00000000000000000000000000000000000000111111111111;
    maze[44] = 50'b00000000000000000000000000000000000000111111111111;
    maze[45] = 50'b11111111111111111111111111111111111111111111111111;
    maze[46] = 50'b11111111111111111111111111111111111111111111111111;
    maze[47] = 50'b11111111111111111111111111111111111111111111111111;
    maze[48] = 50'b11111111111111111111111111111111111111111111111111;
    maze[49] = 50'b11111111111111111111111111111111111111111111111111;


   
    
    
  end
  
endmodule

module alpha2(hpos, vpos, alpha_n);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_n;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-170;
  wire [9:0] y = vpos-200;
  
  assign alpha_n= ((170<=hpos)&(hpos<=219))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
    maze[0]=  50'b110000000000000000000000000000000000000111111111111;
    maze[1]=  50'b111000000000000000000000000000000000000111111111111;
    maze[2]=  50'b111100000000000000000000000000000000000111111111111;
    maze[3]=  50'b111110000000000000000000000000000000000111111111111;
    maze[4]=  50'b111111000000000000000000000000000000000111111111111;
    maze[5]=  50'b111111100000000000000000000000000000000111111111111;
    maze[6]=  50'b111111110000000000000000000000000000000111111111111;
    maze[7]=  50'b111111111000000000000000000000000000000111111111111;
    maze[8]=  50'b111111111100000000000000000000000000000111111111111;
    maze[8]=  50'b111111111110000000000000000000000000000111111111111;
    maze[9]=  50'b111111111111000000000000000000000000000111111111111;
    maze[10]= 50'b111111111111100000000000000000000000000111111111111;
    maze[11]= 50'b111111111111110000000000000000000000000111111111111;
    maze[12]= 50'b111111111111111000000000000000000000000111111111111;
    maze[13]= 50'b111111111111111100000000000000000000000111111111111;
    maze[14]= 50'b111111111111111110000000000000000000000111111111111;
    maze[15]= 50'b111111111111111111000000000000000000000111111111111;
    maze[16]= 50'b111111111111111111100000000000000000000111111111111;
    maze[17]= 50'b111111111111111111110000000000000000000111111111111;
    maze[18]= 50'b111111111111111111111000000000000000000111111111111;
    maze[19]= 50'b111111111111111111111100000000000000000111111111111;
    maze[20]= 50'b111111111111111111111110000000000000000111111111111;
    maze[21]= 50'b111111111111111111111111000000000000000111111111111;
    maze[22]= 50'b111111111111011111111111100000000000000111111111111;
    maze[23]= 50'b111111111111001111111111110000000000000111111111111;
    maze[24]= 50'b111111111111000111111111111000000000000111111111111;
    maze[25]= 50'b111111111111000011111111111100000000000111111111111;
    maze[26]= 50'b111111111111000001111111111110000000000111111111111;
    maze[27]= 50'b111111111111000000111111111111000000000111111111111;
    maze[28]= 50'b111111111111000000011111111111100000000111111111111;

    maze[29]= 50'b111111111111000000001111111111110000000111111111111;

    maze[30]= 50'b111111111111000000000111111111111000000111111111111;
    maze[31]= 50'b111111111111000000000011111111111100000111111111111;
    maze[32]= 50'b111111111111000000000001111111111110000111111111111;
    maze[33]= 50'b111111111111000000000000111111111111000111111111111;
    maze[34]= 50'b111111111111000000000000011111111111100111111111111;
    maze[35]= 50'b111111111111000000000000001111111111110111111111111;
    maze[36]= 50'b111111111111000000000000000111111111111111111111111;
    maze[37]= 50'b111111111111000000000000000011111111111111111111111;
    maze[38]= 50'b111111111111000000000000000001111111111111111111111;
    maze[39]= 50'b111111111111000000000000000000111111111111111111111;

    maze[40]= 50'b111111111111000000000000000000011111111111111111111;
    maze[41]= 50'b111111111111000000000000000000001111111111111111111;
    maze[42]= 50'b111111111111000000000000000000000111111111111111111;
    maze[43]= 50'b111111111111000000000000000000000011111111111111111;
    maze[44]= 50'b111111111111000000000000000000000001111111111111111;
    maze[45]= 50'b111111111111000000000000000000000000111111111111111;
    maze[46]= 50'b111111111111000000000000000000000000011111111111111;
    maze[47]= 50'b111111111111000000000000000000000000001111111111111;
    maze[48]= 50'b111111111111000000000000000000000000000111111111111;
    maze[49]= 50'b111111111111000000000000000000000000000011111111111;
    

   
    
    
  end
  
endmodule
module alpha3(hpos, vpos, alpha_a);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_a;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-250;
  wire [9:0] y = vpos-200;
  
  assign alpha_a= ((250<=hpos)&(hpos<=299))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
    maze[0]  = 50'b11111111111111111111111111111111111111111111111111; 
 	maze[1]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[2]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[3]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[4]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[5]  = 50'b11111111111111111111111111111111111111111111111111;

    maze[6]=  50'b111111111111000000000000000000000000000111111111111;
    maze[7]=  50'b111111111111000000000000000000000000000111111111111;
    maze[8]=  50'b111111111111000000000000000000000000000111111111111;

    maze[8]=  50'b111111111111000000000000000000000000000111111111111;
    maze[9]=  50'b111111111111000000000000000000000000000111111111111;
    maze[10]= 50'b111111111111000000000000000000000000000111111111111;

    maze[11]= 50'b111111111111000000000000000000000000000111111111111;
    maze[12]= 50'b111111111111000000000000000000000000000111111111111;
    maze[13]= 50'b111111111111000000000000000000000000000111111111111;
    maze[14]= 50'b111111111111000000000000000000000000000111111111111;
    maze[15]= 50'b111111111111000000000000000000000000000111111111111;
    maze[16]= 50'b111111111111000000000000000000000000000111111111111;

    maze[17]= 50'b111111111111000000000000000000000000000111111111111;
    maze[18]= 50'b111111111111000000000000000000000000000111111111111;
    maze[19]= 50'b111111111111000000000000000000000000000111111111111;

    maze[20]= 50'b111111111111000000000000000000000000000111111111111;
    maze[21]= 50'b111111111111000000000000000000000000000111111111111;
    maze[22]= 50'b111111111111000000000000000000000000000111111111111;
    maze[23] = 50'b11111111111111111111111111111111111111111111111111;
    maze[24] = 50'b11111111111111111111111111111111111111111111111111;
    maze[25] = 50'b11111111111111111111111111111111111111111111111111;
    maze[26] = 50'b11111111111111111111111111111111111111111111111111;
    maze[27] = 50'b11111111111111111111111111111111111111111111111111;
    maze[28] = 50'b11111111110000000000000000000000000000111111111111;

    maze[29]= 50'b111111111111000000000000000000000000000111111111111;

    maze[30]= 50'b111111111111000000000000000000000000000111111111111;
    maze[31]= 50'b111111111111000000000000000000000000000111111111111;
    maze[32]= 50'b111111111111000000000000000000000000000111111111111;
    maze[33]= 50'b111111111111000000000000000000000000000111111111111;
    maze[34]= 50'b111111111111000000000000000000000000000111111111111;
    maze[35]= 50'b111111111111000000000000000000000000000111111111111;
    maze[36]= 50'b111111111111000000000000000000000000000111111111111;
    maze[37]= 50'b111111111111000000000000000000000000000111111111111;
    maze[38]= 50'b111111111111000000000000000000000000000111111111111;
    maze[39]= 50'b111111111111000000000000000000000000000111111111111;

    maze[40]= 50'b111111111111000000000000000000000000000111111111111;
    maze[41]= 50'b111111111111000000000000000000000000000111111111111;
    maze[42]= 50'b111111111111000000000000000000000000000111111111111;
    maze[43]= 50'b111111111111000000000000000000000000000111111111111;
    maze[44]= 50'b111111111111000000000000000000000000000111111111111;
    maze[45]= 50'b111111111111000000000000000000000000000111111111111;
    maze[46]= 50'b111111111111000000000000000000000000000111111111111;
    maze[47]= 50'b111111111111000000000000000000000000000111111111111;
    maze[48]= 50'b111111111111000000000000000000000000000111111111111;
    maze[49]= 50'b111111111111000000000000000000000000000111111111111;
    

   
    
    
  end
  
endmodule
module alpha5(hpos, vpos, alpha_k);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_k;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-330;
  wire [9:0] y = vpos-200;
  
  assign alpha_k= ((330<=hpos)&(hpos<=379))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
    maze[0]  = 50'b11111111111100000000000000000000000000001111111111;
    maze[1]  = 50'b11111111111100000000000000000000000000011111111110;
    maze[2]  = 50'b11111111111100000000000000000000000000111111111100;
    maze[3]  = 50'b11111111111100000000000000000000000001111111111000;
    maze[4]  = 50'b11111111111100000000000000000000000011111111110000;
    maze[5]  = 50'b11111111111100000000000000000000000111111111100000;
    maze[6]  = 50'b11111111111100000000000000000000001111111111000000;
    maze[7]  = 50'b11111111111100000000000000000000011111111110000000;
    maze[8]  = 50'b11111111111100000000000000000000111111111100000000;
    maze[9]  = 50'b11111111111100000000000000000001111111111000000000;
    maze[10] = 50'b11111111111100000000000000000011111111110000000000;
    maze[11] = 50'b11111111111100000000000000000111111111100000000000;
    maze[12] = 50'b11111111111100000000000000001111111111000000000000;
    maze[13] = 50'b11111111111100000000000000011111111110000000000000;
    maze[14] = 50'b11111111111100000000000000111111111100000000000000;
    maze[15] = 50'b11111111111100000000000001111111111000000000000000;
    maze[16] = 50'b11111111111100000000000011111111110000000000000000;
    maze[17] = 50'b11111111111100000000000111111111100000000000000000;
    maze[18] = 50'b11111111111100000000001111111111000000000000000000;
    maze[19] = 50'b11111111111100000000011111111110000000000000000000;
    maze[20] = 50'b11111111111100000000111111111100000000000000000000;
    maze[21] = 50'b11111111111100000001111111111000000000000000000000;
    maze[22] = 50'b11111111111100000011111111110000000000000000000000;
    maze[23] = 50'b11111111111100000111111111100000000000000000000000;
    maze[24] = 50'b11111111111100001111111111000000000000000000000000;
    maze[25] = 50'b11111111111100011111111110000000000000000000000000;
    maze[26] = 50'b11111111111100111111111100000000000000000000000000;
    maze[27] = 50'b11111111111101111111111000000000000000000000000000;
    maze[28] = 50'b11111111111111111111110000000000000000000000000000;
    maze[29] = 50'b11111111111101111111111000000000000000000000000000;
    maze[30] = 50'b11111111111100111111111100000000000000000000000000;
    maze[31] = 50'b11111111111100011111111110000000000000000000000000;
    maze[32] = 50'b11111111111100001111111111000000000000000000000000;
    maze[33] = 50'b11111111111100000111111111100000000000000000000000;
    maze[34] = 50'b11111111111100000011111111110000000000000000000000;
    maze[35] = 50'b11111111111100000001111111111000000000000000000000;
    maze[36] = 50'b11111111111100000000111111111100000000000000000000;
    maze[37] = 50'b11111111111100000000011111111110000000000000000000;
    maze[38] = 50'b11111111111100000000001111111111000000000000000000;
    maze[39] = 50'b11111111111100000000000111111111100000000000000000;
    maze[40] = 50'b11111111111100000000000011111111110000000000000000;
    maze[41] = 50'b11111111111100000000000001111111111000000000000000;
    maze[42] = 50'b11111111111100000000000000111111111100000000000000;
    maze[43] = 50'b11111111111100000000000000011111111110000000000000;
    maze[44] = 50'b11111111111100000000000000001111111111000000000000;
    maze[45] = 50'b11111111111100000000000000000111111111100000000000;
    maze[46] = 50'b11111111111100000000000000000011111111110000000000;
    maze[47] = 50'b11111111111100000000000000000001111111111000000000;
    maze[48] = 50'b11111111111100000000000000000000111111111100000000;
    maze[49] = 50'b11111111111100000000000000000000011111111110000000;


   
    
    
  end
  
endmodule
module alpha4(hpos, vpos, alpha_e);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_e;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-400;
  wire [9:0] y = vpos-200;
  
  assign alpha_e= ((400<=hpos)&(hpos<=449))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
    maze[0]  = 50'b11111111111111111111111111111111111111111111111111; 
 	maze[1]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[2]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[3]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[4]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[5]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[6]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[7]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[8]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[9]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[10] = 50'b11111111111100000000000000000000000000000000000000;
    maze[11] = 50'b11111111111100000000000000000000000000000000000000;
    maze[12] = 50'b11111111111100000000000000000000000000000000000000;
    maze[13] = 50'b11111111111100000000000000000000000000000000000000;
    maze[14] = 50'b11111111111100000000000000000000000000000000000000;
    maze[15] = 50'b11111111111100000000000000000000000000000000000000;
    maze[16] = 50'b11111111111100000000000000000000000000000000000000;
    maze[17] = 50'b11111111111100000000000000000000000000000000000000;
    maze[18] = 50'b11111111111100000000000000000000000000000000000000;
    maze[19] = 50'b11111111111100000000000000000000000000000000000000;
    maze[20] = 50'b11111111111100000000000000000000000000000000000000;
    maze[21] = 50'b11111111111100000000000000000000000000000000000000;
    maze[22] = 50'b11111111111100000000000000000000000000000000000000;
    maze[23] = 50'b11111111111111111111111111111111111111111111111111;
    maze[24] = 50'b11111111111111111111111111111111111111111111111111;
    maze[25] = 50'b11111111111111111111111111111111111111111111111111;
    maze[26] = 50'b11111111111111111111111111111111111111111111111111;
    maze[27] = 50'b11111111111111111111111111111111111111111111111111;
    maze[28]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[29]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[30]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[31]  = 50'b11111111111100000000000000000000000000000000000000;
    maze[32] = 50'b11111111111100000000000000000000000000000000000000;
    maze[33] = 50'b11111111111100000000000000000000000000000000000000;
    maze[34] = 50'b11111111111100000000000000000000000000000000000000;
    maze[35] = 50'b11111111111100000000000000000000000000000000000000;
    maze[36] = 50'b11111111111100000000000000000000000000000000000000;
    maze[37] = 50'b11111111111100000000000000000000000000000000000000;
    maze[38] = 50'b11111111111100000000000000000000000000000000000000;
    maze[39] = 50'b11111111111100000000000000000000000000000000000000;
    maze[40] = 50'b11111111111100000000000000000000000000000000000000;
    maze[41] = 50'b11111111111100000000000000000000000000000000000000;
    maze[42] = 50'b11111111111100000000000000000000000000000000000000;
    maze[43] = 50'b11111111111100000000000000000000000000000000000000;
    maze[44] = 50'b11111111111100000000000000000000000000000000000000;
    maze[45] = 50'b11111111111111111111111111111111111111111111111111;
    maze[46] = 50'b11111111111111111111111111111111111111111111111111;
    maze[47] = 50'b11111111111111111111111111111111111111111111111111;
    maze[48] = 50'b11111111111111111111111111111111111111111111111111;
    maze[49] = 50'b11111111111111111111111111111111111111111111111111;


   
    
    
  end
  
endmodule
module player1(hpos, vpos, alpha_1);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_1;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-500;
  wire [9:0] y = vpos-200;
  
  assign alpha_1= ((500<=hpos)&(hpos<=549))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
        maze[0]  = 50'b11111111111111111111111111111111111111111111111111; 
 	    maze[1]  = 50'b11111111111111111111111111111111111111111111111111;
        maze[2]  = 50'b11111111111111111111111111111111111111111111111111;
        maze[3]  = 50'b11111111111111111111111111111111111111111111111111;
        maze[4]  = 50'b11111111111111111111111111111111111111111111111111;
        maze[5]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[6] = 50'b00000000000000001111111111111111110000000000000000;
    maze[7] = 50'b00000000000000001111111111111111110000000000000000;
         maze[8]   = 50'b00000000000000001111111111111111110000000000000000;
         maze[9]   = 50'b00000000000000001111111111111111110000000000000000;
         maze[10]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[11]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[12]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[13]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[14]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[15]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[16]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[17]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[18]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[19]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[20]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[21]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[22]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[23]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[24]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[25]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[26]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[27]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[28]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[29]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[30]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[31]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[32]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[33]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[34]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[35]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[36]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[37]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[38]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[39]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[40]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[41]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[42]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[43]  = 50'b00000000000000001111111111111111110000000000000000;
         maze[44]  = 50'b00000000000000001111111111111111110000000000000000;
       
    
    maze[45] = 50'b11111111111111111111111111111111111111111111111111;
    maze[46] = 50'b11111111111111111111111111111111111111111111111111;
    maze[47] = 50'b11111111111111111111111111111111111111111111111111;
    maze[48] = 50'b11111111111111111111111111111111111111111111111111;
    maze[49] = 50'b11111111111111111111111111111111111111111111111111;

    
  end
endmodule

module alpha6(hpos, vpos, alpha_w);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_w;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-200;
  wire [9:0] y = vpos-300;
  
  assign alpha_w= ((200<=hpos)&(hpos<=249))?(((300<=vpos)&(vpos<=349))?maze[y][x]:1'b0):1'b0;
  
  initial begin
    maze[0]= 50'b111111111111000000000000000000000000000111111111111;
    maze[1]= 50'b111111111111000000000000000000000000000111111111111;
    maze[2]= 50'b111111111111000000000000000000000000000111111111111;
    maze[3]= 50'b111111111111000000000000000000000000000111111111111;
    maze[4]=  50'b111111111111000000000000000000000000000111111111111;
    maze[5]=  50'b111111111111000000000000000000000000000111111111111;

    maze[6]=  50'b111111111111000000000000000000000000000111111111111;
    maze[7]=  50'b111111111111000000000000000000000000000111111111111;
    maze[8]=  50'b111111111111000000000000000000000000000111111111111;

    maze[8]=  50'b111111111111000000000000000000000000000111111111111;
    maze[9]=  50'b111111111111000000000000000000000000000111111111111;
    maze[10]= 50'b111111111111000000000000000000000000000111111111111;

    maze[11]= 50'b111111111111000000000000000000000000000111111111111;
    maze[12]= 50'b111111111111000000000000000000000000000111111111111;
    maze[13]= 50'b111111111111000000000000000000000000000111111111111;
    maze[14]= 50'b111111111111000000000000000000000000000111111111111;
    maze[15]= 50'b111111111111000000000000000000000000000111111111111;
    maze[16]= 50'b111111111111000000000000000000000000000111111111111;

    maze[17]= 50'b111111111111000000000000000000000000000111111111111;
    maze[18]= 50'b111111111111000000000000000000000000000111111111111;
    maze[19]= 50'b111111111111000000000000000000000000000111111111111;

    maze[20]= 50'b111111111111000000000000000000000000000111111111111;
    maze[21]= 50'b111111111111000000000000000000000000000111111111111;
    maze[22]= 50'b111111111111000000000000000000000000000111111111111;
    maze[23]= 50'b111111111111000000000000000000000000000111111111111;
    maze[24]= 50'b111111111111000000000000000000000000000111111111111;
    maze[25]= 50'b111111111111000000000000000000000000000111111111111;
    maze[26]= 50'b111111111111000000000000000000000000000111111111111;
    maze[27]= 50'b111111111111000000000000000000000000000111111111111;
    maze[28]= 50'b111111111111000000000000000000000000000111111111111;

    maze[29]= 50'b111111111111000000000000000000000000000111111111111;

    maze[30]= 50'b111111111111000000000111111111000000000111111111111;
    maze[31]= 50'b111111111111000000001111111111100000000111111111111;
    maze[32]= 50'b111111111111000000011111111111110000000111111111111;
    maze[33]= 50'b111111111111000000111111111111111000000111111111111;
    maze[34]= 50'b111111111111000001111111111111111100000111111111111;
    maze[35]= 50'b111111111111000011111111101111111110000111111111111;
    maze[36]= 50'b111111111111000111111111000111111111000111111111111;
    maze[37]= 50'b111111111111111111111110000011111111111111111111111;
    maze[38]= 50'b111111111111111111111100000001111111111111111111111;
    maze[39]= 50'b111111111111111111111000000000111111111111111111111;

    maze[40]= 50'b111111111111111111110000000000011111111111111111111;
    maze[41]= 50'b111111111111111111100000000000001111111111111111111;
    maze[42]= 50'b111111111111111111000000000000000111111111111111111;
    maze[43]= 50'b111111111111111110000000000000000011111111111111111;
    maze[44]= 50'b111111111111111100000000000000000001111111111111111;
    maze[45]= 50'b111111111111111000000000000000000000111111111111111;
    maze[46]= 50'b111111111111110000000000000000000000011111111111111;
    maze[47]= 50'b111111111111100000000000000000000000001111111111111;
    maze[48]= 50'b111111111111000000000000000000000000000111111111111;
    maze[49]= 50'b111111111110000000000000000000000000000011111111111;
    

   
    
    
  end
  
endmodule

module alpha7(hpos, vpos, alpha_o);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_o;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-270;
  wire [9:0] y = vpos-300;
  
  assign alpha_o= ((270<=hpos)&(hpos<=319))?(((300<=vpos)&(vpos<=349))?maze[y][x]:1'b0):1'b0;
  initial begin
    maze[0]= 50'b11111111111111111111111111111111111111111111111111; 
 	maze[1]= 50'b11111111111111111111111111111111111111111111111111;
    maze[2]= 50'b11111111111111111111111111111111111111111111111111;
    maze[3]= 50'b11111111111111111111111111111111111111111111111111;
    maze[4]= 50'b11111111111111111111111111111111111111111111111111;
  maze[5]= 50'b11111111111111111111111111111111111111111111111111;

    maze[6]=  50'b111111111111000000000000000000000000000111111111111;
    maze[7]=  50'b111111111111000000000000000000000000000111111111111;
    maze[8]=  50'b111111111111000000000000000000000000000111111111111;

    maze[8]=  50'b111111111111000000000000000000000000000111111111111;
    maze[9]=  50'b111111111111000000000000000000000000000111111111111;
    maze[10]= 50'b111111111111000000000000000000000000000111111111111;

    maze[11]= 50'b111111111111000000000000000000000000000111111111111;
    maze[12]= 50'b111111111111000000000000000000000000000111111111111;
    maze[13]= 50'b111111111111000000000000000000000000000111111111111;
    maze[14]= 50'b111111111111000000000000000000000000000111111111111;
    maze[15]= 50'b111111111111000000000000000000000000000111111111111;
    maze[16]= 50'b111111111111000000000000000000000000000111111111111;

    maze[17]= 50'b111111111111000000000000000000000000000111111111111;
    maze[18]= 50'b111111111111000000000000000000000000000111111111111;
    maze[19]= 50'b111111111111000000000000000000000000000111111111111;

    maze[20]= 50'b111111111111000000000000000000000000000111111111111;
    maze[21]= 50'b111111111111000000000000000000000000000111111111111;
    maze[22]= 50'b111111111111000000000000000000000000000111111111111;
  maze[23]=  50'b111111111111000000000000000000000000000111111111111;
  maze[24]=  50'b111111111111000000000000000000000000000111111111111;
  maze[25]=  50'b111111111111000000000000000000000000000111111111111;

  maze[26]=  50'b111111111111000000000000000000000000000111111111111;
  maze[27]=  50'b111111111111000000000000000000000000000111111111111;
  maze[28]= 50'b111111111111000000000000000000000000000111111111111;

  maze[29]= 50'b111111111111000000000000000000000000000111111111111;
  maze[30]= 50'b111111111111000000000000000000000000000111111111111;
  maze[31]= 50'b111111111111000000000000000000000000000111111111111;
  maze[32]= 50'b111111111111000000000000000000000000000111111111111;
  maze[33]= 50'b111111111111000000000000000000000000000111111111111;
  maze[34]= 50'b111111111111000000000000000000000000000111111111111;

  maze[35]= 50'b111111111111000000000000000000000000000111111111111;
  maze[36]= 50'b111111111111000000000000000000000000000111111111111;
  maze[37]= 50'b111111111111000000000000000000000000000111111111111;

  maze[38]= 50'b111111111111000000000000000000000000000111111111111;
  maze[39]= 50'b111111111111000000000000000000000000000111111111111;
  maze[40]= 50'b111111111111000000000000000000000000000111111111111;
  maze[41]= 50'b111111111111000000000000000000000000000111111111111;
  maze[42]= 50'b111111111111000000000000000000000000000111111111111;
  maze[43]= 50'b111111111111000000000000000000000000000111111111111;
  
  maze[44] = 50'b11111111111111111111111111111111111111111111111111;
  
  
    maze[45] = 50'b11111111111111111111111111111111111111111111111111;
    maze[46] = 50'b11111111111111111111111111111111111111111111111111;
    maze[47] = 50'b11111111111111111111111111111111111111111111111111;
    maze[48] = 50'b11111111111111111111111111111111111111111111111111;
    maze[49] = 50'b11111111111111111111111111111111111111111111111111;
  
  
  
  
  end
endmodule
module alpha8(hpos, vpos, alpha_n1);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_n1;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-350;
  wire [9:0] y = vpos-300;
  
  assign alpha_n1= ((350<=hpos)&(hpos<=399))?(((300<=vpos)&(vpos<=349))?maze[y][x]:1'b0):1'b0;
  
  initial begin
   maze[0]=  50'b110000000000000000000000000000000000000111111111111;
    maze[1]=  50'b111000000000000000000000000000000000000111111111111;
    maze[2]=  50'b111100000000000000000000000000000000000111111111111;
    maze[3]=  50'b111110000000000000000000000000000000000111111111111;
    maze[4]=  50'b111111000000000000000000000000000000000111111111111;
    maze[5]=  50'b111111100000000000000000000000000000000111111111111;
    maze[6]=  50'b111111110000000000000000000000000000000111111111111;
    maze[7]=  50'b111111111000000000000000000000000000000111111111111;
    maze[8]=  50'b111111111100000000000000000000000000000111111111111;
    maze[8]=  50'b111111111110000000000000000000000000000111111111111;
    maze[9]=  50'b111111111111000000000000000000000000000111111111111;
    maze[10]= 50'b111111111111100000000000000000000000000111111111111;
    maze[11]= 50'b111111111111110000000000000000000000000111111111111;
    maze[12]= 50'b111111111111111000000000000000000000000111111111111;
    maze[13]= 50'b111111111111111100000000000000000000000111111111111;
    maze[14]= 50'b111111111111111110000000000000000000000111111111111;
    maze[15]= 50'b111111111111111111000000000000000000000111111111111;
    maze[16]= 50'b111111111111111111100000000000000000000111111111111;
    maze[17]= 50'b111111111111111111110000000000000000000111111111111;
    maze[18]= 50'b111111111111111111111000000000000000000111111111111;
    maze[19]= 50'b111111111111111111111100000000000000000111111111111;
    maze[20]= 50'b111111111111111111111110000000000000000111111111111;
    maze[21]= 50'b111111111111111111111111000000000000000111111111111;
    maze[22]= 50'b111111111111011111111111100000000000000111111111111;
    maze[23]= 50'b111111111111001111111111110000000000000111111111111;
    maze[24]= 50'b111111111111000111111111111000000000000111111111111;
    maze[25]= 50'b111111111111000011111111111100000000000111111111111;
    maze[26]= 50'b111111111111000001111111111110000000000111111111111;
    maze[27]= 50'b111111111111000000111111111111000000000111111111111;
    maze[28]= 50'b111111111111000000011111111111100000000111111111111;

    maze[29]= 50'b111111111111000000001111111111110000000111111111111;

    maze[30]= 50'b111111111111000000000111111111111000000111111111111;
    maze[31]= 50'b111111111111000000000011111111111100000111111111111;
    maze[32]= 50'b111111111111000000000001111111111110000111111111111;
    maze[33]= 50'b111111111111000000000000111111111111000111111111111;
    maze[34]= 50'b111111111111000000000000011111111111100111111111111;
    maze[35]= 50'b111111111111000000000000001111111111110111111111111;
    maze[36]= 50'b111111111111000000000000000111111111111111111111111;
    maze[37]= 50'b111111111111000000000000000011111111111111111111111;
    maze[38]= 50'b111111111111000000000000000001111111111111111111111;
    maze[39]= 50'b111111111111000000000000000000111111111111111111111;

    maze[40]= 50'b111111111111000000000000000000011111111111111111111;
    maze[41]= 50'b111111111111000000000000000000001111111111111111111;
    maze[42]= 50'b111111111111000000000000000000000111111111111111111;
    maze[43]= 50'b111111111111000000000000000000000011111111111111111;
    maze[44]= 50'b111111111111000000000000000000000001111111111111111;
    maze[45]= 50'b111111111111000000000000000000000000111111111111111;
    maze[46]= 50'b111111111111000000000000000000000000011111111111111;
    maze[47]= 50'b111111111111000000000000000000000000001111111111111;
    maze[48]= 50'b111111111111000000000000000000000000000111111111111;
    maze[49]= 50'b111111111111000000000000000000000000000011111111111;
    

   
    
    
  end
  
endmodule




module player2(hpos, vpos, alpha_2);
  
  input [9:0] hpos;
  input [9:0] vpos;
  output alpha_2;
  
  reg [0:49] maze [0:49];
  
  wire [9:0] x = hpos-500;
  wire [9:0] y = vpos-200;
  
  assign alpha_2= ((500<=hpos)&(hpos<=549))?(((200<=vpos)&(vpos<=249))?maze[y][x]:1'b0):1'b0;
  
  initial begin
         maze[0]  = 50'b11111111111111111111111111111111111111111111111111; 
 	     maze[1]  = 50'b11111111111111111111111111111111111111111111111111;
         maze[2]  = 50'b11111111111111111111111111111111111111111111111111;
         maze[3]  = 50'b11111111111111111111111111111111111111111111111111;
         maze[4]  = 50'b11111111111111111111111111111111111111111111111111;
         maze[5]  = 50'b11111111111111111111111111111111111111111111111111;
    maze[6]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[7]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[8]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[9]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[10]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[11]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[12]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[13]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[14]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[15]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[16]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[17]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[18]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[19]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[20]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[21]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[22]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[23]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[24]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[25]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[26]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[27]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[28]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[29]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[30]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[31]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[32]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[33]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[34]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[35]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[36]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[37]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[38]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[39]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[40]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[41]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[41]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[42]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[43]  =       50'b0000000000011111111111100000111111111110000000000;
    maze[44]  =       50'b0000000000011111111111100000111111111110000000000;

    
         maze[45] = 50'b11111111111111111111111111111111111111111111111111;
         maze[46] = 50'b11111111111111111111111111111111111111111111111111;
         maze[47] = 50'b11111111111111111111111111111111111111111111111111;
         maze[48] = 50'b11111111111111111111111111111111111111111111111111;
         maze[49] = 50'b11111111111111111111111111111111111111111111111111;

    
  end
endmodule

module snaketop(
  input clk_d,
  input clk_u,
  input reg [4:0] state_snake1,
  input reg [4:0] state_snake2,
  input [9:0] x, 
  input [9:0] y,
  input video_on,
  output reg [3:0] red,
  output reg [3:0] green ,
  output reg [3:0] blue );
  
 reg reset=0;
  
  reg square; 
  reg snake;
  reg snake1, snake2, snake3, snake4;
  reg food;
  reg foodeat = 0;
  
  //snake 2
  reg snake2_head; //head of the snake
  reg snake2_1, snake2_2, snake2_3, snake2_4;
  //
  
  reg [9:0] headx=200;
  reg [8:0] heady = 150;
  reg [9:0] headx1 = 200;
  reg [8:0] heady1 = 130;
  reg [9:0] headx2 = 200;
  reg [8:0] heady2 = 110;
  reg [9:0] headx3 = 220;
  reg [8:0] heady3= 110;
  reg [9:0] headx4 = 240;
  reg [8:0] heady4 = 110;
  
  reg [9:0] foodx = 300;
  reg [8:0] foody = 200;
  
  reg [2:0] gs_S1, gs_S2, ns_S1, ns_S2;
  
  //snake 2
  reg [9:0] head2_x=560;
  reg [8:0] head2_y = 100;
  reg [9:0] head2_x1 = 560;
  reg [8:0] head2_y1 = 80;
  reg [9:0] head2_x2 = 560;
  reg [8:0] head2_y2 = 60;
  reg [9:0] head2_x3 = 580;
  reg [8:0] head2_y3= 60;
  reg [9:0] head2_x4 = 600;
  reg [8:0] head2_y4 = 60;
 
  //reg [4:0] dir2;
  
//  always@(posedge clk_d)
//    begin 
//    if (R) 
//    dir2 = 5'b10001;
//    if (D)
//    dir2 = 5'b11010;
//    if (L) 
//    dir2 = 5'b00101;
//    if (U)
//    dir2 = 5'b10101;
//    end 
  
  reg food_collide_S1, food_collide_S2;
  reg bCollision_1, bCollision_2;

reg snake1_score, snake2_score;
reg [9:0] s1s1x, s1s2x, s1s3x, s1s4x, s2s1x, s2s2x, s2s3x, s2s4x;
reg [8:0] s1s1y, s1s2y, s1s3y, s1s4y, s2s1y, s2s2y, s2s3y, s2s4y;
      
//reg [9:0] s1s1x=0, s1s2x=0, s1s3x=0, s1s4x=0, s2s1x=0, s2s2x=0, s2s3x=0, s2s4x=0;
//reg [8:0] s1s1y=0, s1s2y=0, s1s3y=0, s1s4y=0, s2s1y=0, s2s2y=0, s2s3y=0, s2s4y=0;
      
  
  parameter START = 3'b000; 
  parameter One_Point = 3'b001; 
  parameter Two_Points = 3'b010;
  parameter Three_Points = 3'b011;
  parameter Four_Points = 3'b100;
  parameter WON = 3'b101;
  parameter LOST = 3'b110;

  wire alpha_S;
  wire alpha_N;
  wire alpha_A;
  
  wire alpha_E;
  wire alpha_K;
  wire alpha_1;
  wire alpha_2;
  wire alpha_W;
  wire alpha_O;
  wire alpha_N1;


alpha1 a1( .hpos(x),
          .vpos(y),
  .alpha_s(alpha_S));
  
alpha2 a2( .hpos(x),
  .vpos(y),
   .alpha_n(alpha_N));
  
   alpha3 a3( .hpos(x),
  .vpos(y),
   .alpha_a(alpha_A));
  
  
   alpha4 a4( .hpos(x),
  .vpos(y),
   .alpha_e(alpha_E));
  
   alpha5 a5( .hpos(x),
  .vpos(y),
   .alpha_k(alpha_K));
  
   alpha6 a6( .hpos(x),
  .vpos(y),
   .alpha_w(alpha_W));
  
   alpha7 a7( .hpos(x),
  .vpos(y),
   .alpha_o(alpha_O));
  
   alpha8 a8( .hpos(x),
  .vpos(y),
    .alpha_n1(alpha_N1));
  
  
  player1 p1( .hpos(x),
  .vpos(y),
    .alpha_1(alpha_1));

  player2 p2( .hpos(x),
  .vpos(y),
  .alpha_2(alpha_2));
  
  initial gs_S1 = START;
initial gs_S2 = START;

  //reg reset=0;
  
//   if (state_snake1 == 5'b11111)
//       begin 
////            headx <= 20;
////            heady <= 20;
//            reset =1;
//       end
 
 
 
  //always @ (posedge clk_u or posedge reset) 
  always@(posedge clk_u)
  begin
    


food_collide_S1 = (((headx - foodx < 20) & (headx - foodx > 0)) || ((foodx - headx > 0) & (foodx - headx < 20))) & (((heady - foody < 20) & (heady - foody > 0)) || ((foody - heady < 20)) & (foody - heady > 0));
    
    
food_collide_S2 = (((head2_x - foodx < 20) & (head2_x - foodx > 0)) || ((foodx - head2_x > 0) & (foodx - head2_x < 20))) & (((head2_y - foody < 20) & (head2_y - foody > 0)) || ((foody - head2_y < 20)) & (foody - head2_y > 0));
    
    
    if (food_collide_S1 || food_collide_S2)
      foodeat = 1;
    
    
bCollision_1 =  (((((headx - head2_x1  < 20) & (headx - head2_x1  > 0)) || ((head2_x1  - headx > 0) & (head2_x1  - headx < 20))) & (((heady - head2_y1 < 20) & (heady - head2_y1> 0)) || ((head2_y1- heady < 20)) & (head2_y1 - heady > 0))) || ((((headx - head2_x2  < 20) & (headx - head2_x2  > 0)) || ((head2_x2  - headx > 0) & (head2_x2  - headx < 20))) & (((heady - head2_y2 < 20) & (heady - head2_y2 > 0)) || ((head2_y2- heady < 20)) & (head2_y2 - heady > 0))) || ((((headx - head2_x3  < 20) & (headx - head2_x3  > 0)) || ((head2_x3  - headx > 0) & (head2_x3  - headx < 20))) & (((heady - head2_y3 < 20) & (heady - head2_y3> 0)) || ((head2_y3- heady < 20)) & (head2_y3 - heady > 0))) || ((((headx - head2_x4  < 20) & (headx - head2_x4  > 0)) || ((head2_x4  - headx > 0) & (head2_x4  - headx < 20))) & (((heady - head2_y4 < 20) & (heady - head2_y4> 0)) || ((head2_y4- heady < 20)) & (head2_y4 - heady > 0))));
    

bCollision_2 = (((((head2_x - headx1 < 20) & (head2_x - headx1 > 0)) || ((headx1 - head2_x > 0) & (headx1 - head2_x < 20))) & (((head2_y - heady1 < 20) & (head2_y - heady1 > 0)) || ((heady1- head2_y < 20)) & (heady1 - head2_y > 0))) || ((((head2_x - headx2 < 20) & (head2_x - headx2 > 0)) || ((headx2 - head2_x > 0) & (headx2 - head2_x < 20))) & (((head2_y- heady2 < 20) & (head2_y - heady2 > 0)) || ((heady2- head2_y < 20)) & (heady2 - head2_y > 0))) || ((((head2_x - headx3 < 20) & (head2_x- headx3 > 0)) || ((headx3 - head2_x > 0) & (headx3 - head2_x< 20))) & (((head2_y - heady3 < 20) & (head2_y- heady3 > 0)) || ((heady3- head2_y < 20)) & (heady3 - head2_y > 0))) || ((((head2_x - headx4 < 20) & (head2_x- headx4 > 0)) || ((headx4 - head2_x > 0) & (headx4 - head2_x< 20))) & (((head2_y - heady4 < 20) & (head2_y- heady4 > 0)) || ((heady4 - head2_y < 20)) & (heady4 - head2_y > 0))));  
    
    if (state_snake1 == 5'b11111)
            reset =1;

  	case (gs_S1)
    START:
      begin
      if (food_collide_S1)
        ns_S1 = One_Point;
      else if (bCollision_1)
        ns_S1 = LOST;
      else 
        ns_S1 = START;
      end
    One_Point:
      begin
      if (food_collide_S1)
        ns_S1 = Two_Points;
      else if (bCollision_1)
        ns_S1 = LOST;
      else 
        ns_S1 = One_Point;
      end
    Two_Points:
      begin
      if (food_collide_S1)
        ns_S1 = Three_Points;
      else if (bCollision_1)
        ns_S1 = LOST;
      else 
        ns_S1 = Two_Points;
      end
    Three_Points:
      begin
      if (food_collide_S1)
        ns_S1 = Four_Points;
      else if (bCollision_1)
        ns_S1 = LOST;
      else 
        ns_S1 = Three_Points;
      end
    Four_Points:
      begin
      if (food_collide_S1)
        ns_S1 = WON;
      else if (bCollision_1)
        ns_S1 = LOST;
      else 
        ns_S1 = Four_Points;
      end
    WON:
      begin
        ns_S1 = WON;
      end
    LOST:
      begin
        ns_S1 = LOST;
       end
    default:
      ns_S1 = START;
  endcase
  gs_S1 = ns_S1;
        
        
        
  case (gs_S2)
    START:
      begin
     if (food_collide_S2)
        ns_S2 = One_Point;
     else if (bCollision_2)
        ns_S2 = LOST;
      else 
        ns_S2 = START;
      end
    One_Point:
      begin
      if (food_collide_S2)
        ns_S2 = Two_Points;
      else if (bCollision_2)
        ns_S2 = LOST;
      else 
        ns_S2 = One_Point;
      end
    Two_Points:
      begin
      if (food_collide_S2)
        ns_S2 = Three_Points;
      else if (bCollision_2)
        ns_S2 = LOST;
      else 
        ns_S2 = Two_Points;
      end
    Three_Points:
      begin
      if (food_collide_S2)
        ns_S2 = Four_Points;
      else if (bCollision_1)
        ns_S2 = LOST;
      else 
        ns_S2 = Three_Points;
      end
    Four_Points:
      begin
      if (food_collide_S2)
        ns_S2 = WON;
      else if (bCollision_2)
        ns_S2 = LOST;
      else 
        ns_S2 = Four_Points;
      end
    WON:
        begin
        ns_S2 = WON;
        end
        
    LOST:
        begin
        ns_S2 = LOST;
      
        end
    default:
      ns_S2 = START;
  endcase
    

  gs_S2 = ns_S2;
        
        
        if (reset==1)
        begin
        gs_S1 = START;
        gs_S2 = START;
        end
  
  	
    
    if (foodeat)
        begin 
         foodx = 80 + (headx *2 + headx1*2 + headx2) % 450;
         foody = 80 + (heady*2 + headx1) %320;
         foodeat = 0;
         food_collide_S1 = 0;
          food_collide_S2 = 0;
        end 
         

       
       heady1 <= heady; 
       headx1 <= headx;
       heady2 <= heady1;
       headx2 <= headx1;
       heady3 <= heady2;
       headx3 <= headx2;
       heady4 <= heady3;
       headx4 <= headx3;
      
       
//      if (dir == 5'b00100)
//        headx <= headx - 15;
//      else if (dir == 5'b00010)
//        heady <= heady - 15;
//      else if (dir == 5'b01000)
//        heady <= heady + 15;
//      else if (dir == 5'b10000)
//        headx <= headx + 15;
        
         if (state_snake1 == 5'b00100)
        headx <= headx - 15;
      else if (state_snake1 == 5'b00010)
        heady <= heady - 15;
      else if (state_snake1 == 5'b01000)
        heady <= heady + 15;
      else if (state_snake1 == 5'b10000)
        headx <= headx + 15;
      else if (state_snake1 == 5'b11111)
       begin 
//            headx <= 20;
//            heady <= 20;
            reset =1;
       end
 
 
  
       head2_y1 <= head2_y; 
       head2_x1 <= head2_x;
       head2_y2 <= head2_y1;
       head2_x2 <= head2_x1;
       head2_y3 <= head2_y2;
       head2_x3 <= head2_x2;
       head2_y4 <= head2_y3;
       head2_x4 <= head2_x3;
       
//       if (state_snake2== 5'b00100)
//        head2_x <= head2_x - 15;
//      else if (state_snake2 == 5'b00010)
//        head2_y <= head2_y - 15;
//      else if (state_snake2 == 5'b01000)
//        head2_y <= head2_y + 15;
//      else if (state_snake2 == 5'b10001)
//        head2_x <= head2_x + 15;
        
        if (state_snake2 == 5'b00100)
        head2_x <= head2_x - 15;
      else if (state_snake2 == 5'b00010)
        head2_y <= head2_y - 15;
      else if (state_snake2 == 5'b01000)
        head2_y <= head2_y + 15;
      else if (state_snake2 == 5'b10000)
        head2_x <= head2_x + 15;
   if ((gs_S1 == START)  && (gs_S2 == START))
        begin
        //snake1_score=0; snake2_score=0;
s1s1x=0; s1s2x=0; s1s3x=0; s1s4x=0; s2s1x=0; s2s2x=0; s2s3x=0; s2s4x=0;
s1s1y=0; s1s2y=0; s1s3y=0; s1s4y=0; s2s1y=0; s2s2y=0; s2s3y=0; s2s4y=0;
        end
   if (gs_S1 == One_Point)
        begin
          s1s1x = 20;
          s1s1y = 20;
        end
      if (gs_S1 == Two_Points)
        begin
          s1s2x = 30;
          s1s2y = 20;
        end
      if (gs_S1 == Three_Points)
        begin
          s1s3x = 40;
          s1s3y = 20;
        end
      if (gs_S1 == Four_Points)
        begin
          s1s4x = 50;
          s1s4y = 20;
        end
      
      
      if (gs_S2 == One_Point)
        begin
          s2s1x = 600;
          s2s1y = 20;
        end
      if (gs_S2 == Two_Points)
        begin
          s2s2x = 590;
          s2s2y = 20;
        end
      if (gs_S2 == Three_Points)
        begin
          s2s3x = 580;
          s2s3y = 20;
        end
      if (gs_S2 == Four_Points)
        begin
          s2s4x = 570;
          s2s4y = 20;
        end
         
   end

   
   
   
       

 
  //always @(posedge clk_d or posedge reset)
  always @(posedge clk_d )
  begin
      
    square = (x>0) & (x<620) & (y>0) & (y< 460);
    snake = (x > headx) & (x < headx + 20) & (y>heady) & (y<heady + 20); 
    snake1 = (x > headx1) & (x < headx1 + 20) & (y>heady1) & (y<heady1 + 20);
    snake2 = (x > headx2) & (x < headx2 + 20) & (y>heady2) & (y<heady2 + 20);
    snake3 = (x > headx3) & (x < headx3 + 20) & (y>heady3) & (y<heady3 + 20);
    snake4 = (x > headx4) & (x < headx4 + 20) & (y>heady4) & (y<heady4 + 20);
    
    //snake 2
     
     snake2_head = (x > head2_x) & (x < head2_x + 20) & (y > head2_y) & (y<head2_y +20);
     snake2_1 = (x > head2_x1)& (x < head2_x1+ 20) & (y > head2_y1) & (y<head2_y1+20);
     snake2_2= (x > head2_x2)& (x < head2_x2+ 20) & (y > head2_y2) & (y<head2_y2+20);
     snake2_3 = (x > head2_x3)& (x < head2_x3+ 20) & (y > head2_y3) & (y<head2_y3+20);
     snake2_4 = (x > head2_x4)& (x < head2_x4+ 20) & (y > head2_y4) & (y<head2_y4+20);
     //
    
    food = (x > foodx) & (x < foodx + 20) & (y> foody) & (y<foody + 20); 
    
    snake1_score = (((x > s1s1x) & (x < s1s1x + 5) & (y> s1s1y) & (y< s1s1y + 5)) || ((x > s1s2x) & (x < s1s2x + 5) & (y> s1s2y) & (y< s1s2y + 5)) || ((x > s1s3x) & (x < s1s3x + 5) & (y> s1s3y) & (y< s1s3y + 5)) || ((x > s1s4x) & (x < s1s4x + 5) & (y> s1s4y) & (y< s1s4y + 5)));
      
    snake2_score = (((x > s2s1x) & (x < s2s1x + 5) & (y> s2s1y) & (y< s2s1y + 5)) || ((x > s2s2x) & (x < s2s2x + 5) & (y> s2s2y) & (y< s2s2y + 5)) || ((x > s2s3x) & (x < s2s3x + 5) & (y> s2s3y) & (y< s2s3y + 5)) || ((x > s2s4x) & (x < s2s4x + 5) & (y> s2s4y) & (y< s2s4y + 5)));
    end
    
  
  //always @ (posedge clk_d or posedge reset) 
  always @ (posedge clk_d ) 
    begin 
      if ((gs_S1 == WON) || (gs_S2 == LOST))
        begin 
           red <= 4'h0;
    green <=(alpha_S||alpha_N||alpha_A||alpha_K||alpha_E||alpha_1||alpha_W||alpha_O||alpha_N1)? 4'hF:4'h0;
    blue<=(alpha_S||alpha_N||alpha_A||alpha_K||alpha_E||alpha_1||alpha_W||alpha_O||alpha_N1)? 4'hF:4'h0;
        reset=0;
        end
      
      else if ((gs_S2 == WON) || (gs_S1 == LOST))
        begin 
           red <=  (alpha_S||alpha_N||alpha_A||alpha_K||alpha_E||alpha_2||alpha_W||alpha_O||alpha_N1)? 4'hF:4'h0;
    green <=  (alpha_S||alpha_N||alpha_A||alpha_K||alpha_E||alpha_2||alpha_W||alpha_O||alpha_N1)? 4'hF:4'h0;
    blue<=4'h0;
        reset=0;
        end
        
      else 
        begin
        
//      green[1] = ~(snake||food|| snake1|| snake2 || snake3 || snake4 || snake2_head||snake2_1|| snake2_2|| snake2_3|| snake2_4);
//      blue[1] = (snake||food|| snake1|| snake2 || snake3 || snake4) ;
//      red[3] = (food || snake2_head||snake2_1|| snake2_2|| snake2_3|| snake2_4);
red <= (food || snake2_head||snake2_1|| snake2_2|| snake2_3|| snake2_4)? 4'hF:4'h0;
blue <= (snake||food|| snake1|| snake2 || snake3 || snake4)? 4'hF:4'h0;
green = (snake1_score || snake2_score)? 4'hF: 4'h0;
        end
    end
 
endmodule
